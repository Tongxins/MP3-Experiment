library verilog;
use verilog.vl_types.all;
entity eight2deightconcat_sv_unit is
end eight2deightconcat_sv_unit;
