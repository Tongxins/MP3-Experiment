library verilog;
use verilog.vl_types.all;
entity sixteen2donetwentyeightconcat_sv_unit is
end sixteen2donetwentyeightconcat_sv_unit;
