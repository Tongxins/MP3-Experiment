library verilog;
use verilog.vl_types.all;
entity zextlshf_sv_unit is
end zextlshf_sv_unit;
