library verilog;
use verilog.vl_types.all;
entity bytefill_sv_unit is
end bytefill_sv_unit;
