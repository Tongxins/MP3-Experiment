library verilog;
use verilog.vl_types.all;
entity l1dcache_control_sv_unit is
end l1dcache_control_sv_unit;
