library verilog;
use verilog.vl_types.all;
entity l1icache_sv_unit is
end l1icache_sv_unit;
