library verilog;
use verilog.vl_types.all;
entity lshf1_sv_unit is
end lshf1_sv_unit;
