library verilog;
use verilog.vl_types.all;
entity shft_sv_unit is
end shft_sv_unit;
