library verilog;
use verilog.vl_types.all;
entity sixteenbitadder_sv_unit is
end sixteenbitadder_sv_unit;
