library verilog;
use verilog.vl_types.all;
entity hazardDetection_sv_unit is
end hazardDetection_sv_unit;
