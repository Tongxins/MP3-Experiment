library verilog;
use verilog.vl_types.all;
entity csreg_sv_unit is
end csreg_sv_unit;
