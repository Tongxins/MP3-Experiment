library verilog;
use verilog.vl_types.all;
entity l2cache_datapath_sv_unit is
end l2cache_datapath_sv_unit;
