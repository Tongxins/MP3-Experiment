library verilog;
use verilog.vl_types.all;
entity l1cache_datapath_sv_unit is
end l1cache_datapath_sv_unit;
