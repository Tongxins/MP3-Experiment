library verilog;
use verilog.vl_types.all;
entity l2cache_control_sv_unit is
end l2cache_control_sv_unit;
